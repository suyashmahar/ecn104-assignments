 module module_name( ...module_input_and_outputs... );
   ...
   // Module functionality
   ...
 endmodule; 
