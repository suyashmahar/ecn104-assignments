...
  always @( ...condition... ) begin
      ...
      // Description of conditional event
      ...
  end
...
   
