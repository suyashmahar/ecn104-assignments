`timescale 1ns/1ps

module module_1_1_ (input [31:0] inputSignal, output [31:0] result);
    assign result = inputSignal << 5;
endmodule
