  module andGate (inputA, inputB, result);
         ...
         // AND gate functionality
         ...
  endmodule
